`timescale 1ns/1ps
module sr_flip_flop (
    input S,
    input R,
    input clk,
    input reset,
    output reg Q,
    output reg Qn
);

always @(posedge clk or posedge reset) begin
    if (reset) begin
        Q <= 0;
        Qn <= 1;
    end else begin
        case ({S, R})
            2'b00: ;            // No change
            2'b01: begin        // Reset
                Q <= 0;
                Qn <= 1;
            end
            2'b10: begin        // Set
                Q <= 1;
                Qn <= 0;
            end
            2'b11: begin        
                Q <= 1'bx;
                Qn <= 1'bx;
            end
        endcase
    end
end

endmodule
