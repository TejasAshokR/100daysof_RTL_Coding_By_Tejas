`timescale 1ns/1ps
module test_bench;
reg [2:0]i;
wire [7:0]out;
decoder dut(i,out);
initial
begin
i=3'b000;
#10;
end
always begin
      #10 i=3'b000;
	   #10 i=3'b001;
		#10 i=3'b010;
	   #10 i=3'b011;
	   #10 i=3'b100;
	   #10 i=3'b101;
		#10 i=3'b110;
		#10 i=3'b111;
end
initial begin
$monitor("i=%b out=%b",i,out);
#90 $finish;
end
endmodule
